CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
90 0 2 120 10
176 83 1278 749
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 179 457 276
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 941 177 0 1 11
0 12
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
40346 0
0
2 +V
167 940 318 0 1 3
0 4
0
0 0 53728 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6957 0 0
2
40346 1
0
7 Ground~
168 939 350 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8646 0 0
2
40346 2
0
7 Pulser~
4 940 414 0 10 12
0 28 29 5 30 0 0 10 10 9
8
0
0 0 4128 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3721 0 0
2
40346 3
0
14 Logic Display~
6 1407 118 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
436 0 0
2
40346 4
0
6 74LS95
110 1375 255 0 12 25
0 12 5 5 4 2 11 10 9 7
31 32 33
0
0 0 4320 0
6 74LS95
-21 -51 21 -43
3 U11
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
6694 0 0
2
40346 5
0
6 74LS95
110 1217 254 0 12 25
0 12 5 5 6 3 4 4 8 9
34 35 36
0
0 0 4320 0
6 74LS95
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
6682 0 0
2
40346 6
0
6 74LS95
110 1058 254 0 12 25
0 12 5 5 2 2 4 4 4 8
37 38 39
0
0 0 4320 0
6 74LS95
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
5326 0 0
2
40346 7
0
2 +V
167 84 437 0 1 3
0 13
0
0 0 53728 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7444 0 0
2
5.89481e-315 0
0
10 2-In NAND~
219 764 249 0 3 22
0 10 6 21
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 8 0
1 U
364 0 0
2
5.89481e-315 5.26354e-315
0
10 2-In NAND~
219 765 337 0 3 22
0 10 19 20
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
3314 0 0
2
5.89481e-315 5.30499e-315
0
10 2-In NAND~
219 574 229 0 3 22
0 18 17 16
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
5933 0 0
2
5.89481e-315 5.32571e-315
0
10 2-In NAND~
219 523 202 0 3 22
0 6 15 18
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 7 0
1 U
9123 0 0
2
5.89481e-315 5.34643e-315
0
10 2-In NAND~
219 523 258 0 3 22
0 11 3 17
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
3297 0 0
2
5.89481e-315 5.3568e-315
0
10 2-In NAND~
219 333 249 0 3 22
0 23 15 22
0
0 0 96 0
6 74LS00
-14 -24 28 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 82
65 0 0 0 4 2 7 0
1 U
3530 0 0
2
5.89481e-315 5.36716e-315
0
10 2-In NAND~
219 124 153 0 3 22
0 26 25 24
0
0 0 96 512
6 74LS00
-14 -24 28 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 26
65 0 0 0 4 1 7 0
1 U
7522 0 0
2
5.89481e-315 5.37752e-315
0
6 JK RN~
219 651 266 0 6 22
0 16 14 11 13 23 10
0
0 0 4448 0
2 01
-8 -42 6 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 3 0
1 U
5284 0 0
2
40346 8
0
10 3-In NAND~
219 194 174 0 4 22
0 6 10 11 25
0
0 0 96 180
6 74LS10
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 4 0
1 U
3779 0 0
2
40346 9
0
10 3-In NAND~
219 195 133 0 4 22
0 19 23 15 26
0
0 0 96 180
6 74LS10
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 118
65 0 0 0 3 1 4 0
1 U
4727 0 0
2
40346 10
0
7 Pulser~
4 83 372 0 10 12
0 40 41 14 42 0 0 10 10 9
8
0
0 0 4128 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3907 0 0
2
5.89481e-315 5.38788e-315
0
14 Logic Display~
6 605 60 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4934 0 0
2
5.89481e-315 5.39306e-315
0
14 Logic Display~
6 560 60 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3945 0 0
2
5.89481e-315 5.39824e-315
0
14 Logic Display~
6 514 60 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7226 0 0
2
5.89481e-315 5.40342e-315
0
14 Logic Display~
6 467 60 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3492 0 0
2
5.89481e-315 5.4086e-315
0
6 JK RN~
219 860 266 0 6 22
0 21 14 20 13 15 11
0
0 0 4448 0
2 00
-8 -42 6 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 2 0
1 U
366 0 0
2
40346 11
0
6 JK RN~
219 417 266 0 6 22
0 22 14 13 13 19 6
0
0 0 4448 0
2 02
-8 -42 6 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 20729136
65 0 0 0 2 2 1 0
1 U
3477 0 0
2
40346 12
0
6 JK RN~
219 205 266 0 6 22
0 24 14 13 13 43 3
0
0 0 4448 0
2 03
-8 -42 6 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 20730052
65 0 0 512 2 1 1 0
1 U
3299 0 0
2
40346 13
0
65
5 0 3 0 0 12416 0 7 0 0 51 4
1185 263
1167 263
1167 83
467 83
8 0 4 0 0 4096 0 8 0 0 6 2
1026 290
1002 290
3 0 5 0 0 4096 0 6 0 0 4 2
1337 246
1286 246
0 2 5 0 0 8192 0 0 6 23 0 4
1132 405
1286 405
1286 237
1337 237
7 0 4 0 0 0 0 8 0 0 6 2
1026 281
1002 281
6 0 4 0 0 8192 0 8 0 0 18 3
1026 272
1002 272
1002 327
7 0 4 0 0 0 0 7 0 0 8 2
1185 281
1167 281
6 0 4 0 0 0 0 7 0 0 18 3
1185 272
1167 272
1167 327
5 0 2 0 0 4096 0 8 0 0 10 2
1026 263
1016 263
4 0 2 0 0 8192 0 8 0 0 17 3
1026 254
1016 254
1016 344
4 0 6 0 0 12416 0 7 0 0 50 4
1185 254
1177 254
1177 93
514 93
9 1 7 0 0 4224 0 6 5 0 0 2
1407 264
1407 136
8 9 8 0 0 4224 0 7 8 0 0 4
1185 290
1121 290
1121 263
1090 263
8 9 9 0 0 4224 0 6 7 0 0 4
1343 291
1274 291
1274 263
1249 263
7 0 10 0 0 12416 0 6 0 0 49 4
1343 282
1328 282
1328 103
560 103
6 0 11 0 0 12416 0 6 0 0 48 4
1343 273
1317 273
1317 114
605 114
1 5 2 0 0 4224 0 3 6 0 0 4
939 344
1307 344
1307 264
1343 264
4 1 4 0 0 12416 0 6 2 0 0 4
1343 255
1297 255
1297 327
940 327
1 0 12 0 0 8192 0 6 0 0 20 3
1343 228
1343 177
1185 177
1 0 12 0 0 8320 0 7 0 0 21 3
1185 227
1185 177
1026 177
1 1 12 0 0 0 0 8 1 0 0 3
1026 227
1026 177
953 177
3 0 5 0 0 0 0 7 0 0 23 2
1179 245
1132 245
2 0 5 0 0 8320 0 7 0 0 25 4
1179 236
1132 236
1132 405
989 405
3 0 5 0 0 0 0 8 0 0 25 2
1020 245
989 245
2 3 5 0 0 0 0 8 4 0 0 4
1020 236
989 236
989 405
964 405
3 0 13 0 0 4096 0 26 0 0 30 3
393 267
393 306
417 306
3 0 13 0 0 0 0 27 0 0 31 3
181 267
181 306
205 306
0 4 13 0 0 4096 0 0 25 29 0 3
651 446
860 446
860 297
4 0 13 0 0 8320 0 17 0 0 30 3
651 297
651 446
417 446
4 0 13 0 0 0 0 26 0 0 31 3
417 297
417 446
205 446
1 4 13 0 0 0 0 9 27 0 0 3
84 446
205 446
205 297
0 2 14 0 0 4096 0 0 25 33 0 4
605 363
824 363
824 258
829 258
0 2 14 0 0 4224 0 0 17 34 0 4
386 363
606 363
606 258
620 258
0 2 14 0 0 0 0 0 26 35 0 3
174 363
386 363
386 258
2 3 14 0 0 0 0 27 20 0 0 3
174 258
174 363
107 363
1 0 11 0 0 0 0 14 0 0 61 3
499 249
488 249
488 165
2 0 15 0 0 4096 0 13 0 0 60 2
499 211
499 124
3 1 16 0 0 12416 0 12 17 0 0 4
601 229
606 229
606 249
627 249
6 2 3 0 0 0 0 27 14 0 0 6
229 249
262 249
262 323
487 323
487 267
499 267
1 0 6 0 0 0 0 13 0 0 65 2
499 193
441 193
3 2 17 0 0 4224 0 14 12 0 0 2
550 258
550 238
3 1 18 0 0 4224 0 13 12 0 0 2
550 202
550 220
2 6 6 0 0 0 0 10 26 0 0 6
740 258
702 258
702 297
470 297
470 249
441 249
1 0 10 0 0 0 0 10 0 0 46 4
740 240
726 240
726 249
690 249
2 5 19 0 0 12288 0 11 26 0 0 6
741 346
678 346
678 311
461 311
461 267
447 267
1 6 10 0 0 0 0 11 17 0 0 4
741 328
690 328
690 249
675 249
3 0 11 0 0 0 0 17 0 0 61 3
627 267
617 267
617 165
1 0 11 0 0 0 0 21 0 0 61 2
605 78
605 165
1 0 10 0 0 0 0 22 0 0 63 2
560 78
560 174
0 1 6 0 0 0 0 0 23 65 0 4
422 183
422 100
514 100
514 78
6 1 3 0 0 0 0 27 24 0 0 4
229 249
229 90
467 90
467 78
3 3 20 0 0 8320 0 11 25 0 0 4
792 337
793 337
793 267
836 267
3 1 21 0 0 4224 0 10 25 0 0 2
791 249
836 249
1 3 22 0 0 4224 0 26 15 0 0 2
393 249
360 249
0 2 15 0 0 4096 0 0 15 60 0 3
278 124
278 258
309 258
0 1 23 0 0 4096 0 0 15 62 0 3
290 133
290 240
309 240
3 1 24 0 0 8320 0 16 27 0 0 4
99 153
98 153
98 249
181 249
4 2 25 0 0 8320 0 18 16 0 0 4
167 174
158 174
158 162
150 162
4 1 26 0 0 8320 0 19 16 0 0 4
168 133
158 133
158 144
150 144
5 3 15 0 0 8320 0 25 19 0 0 3
890 267
890 124
219 124
6 3 11 0 0 0 0 25 18 0 0 3
884 249
884 165
218 165
5 2 23 0 0 8320 0 17 19 0 0 3
681 267
681 133
219 133
6 2 10 0 0 0 0 17 18 0 0 3
675 249
675 174
218 174
5 1 19 0 0 8320 0 26 19 0 0 3
447 267
447 142
219 142
6 1 6 0 0 0 0 26 18 0 0 3
441 249
441 183
218 183
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
