CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
370 0 2 80 10
176 83 1278 749
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 179 457 276
9437202 0
0
6 Title:
5 Name:
0
0
0
34
2 +V
167 940 318 0 1 3
0 6
0
0 0 53744 0
2 5V
-8 -22 6 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4518 0 0
2
5.8948e-315 0
0
7 Ground~
168 939 350 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7215 0 0
2
5.8948e-315 0
0
7 Pulser~
4 940 414 0 10 12
0 32 33 7 34 0 0 1 1 1
8
0
0 0 4144 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3532 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1407 118 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6722 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1275 468 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7596 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1296 468 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 LSB
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5232 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1254 468 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7795 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1232 469 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6312 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1181 469 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8435 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1159 469 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3561 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1137 469 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 C6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9517 0 0
2
5.8948e-315 0
0
14 Logic Display~
6 1114 469 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 MSB
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3167 0 0
2
5.8948e-315 0
0
6 74LS95
110 1375 255 0 12 25
0 18 7 7 6 2 17 16 8 15
35 3 4
0
0 0 4336 0
6 74LS95
-21 -51 21 -43
3 U11
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
3315 0 0
2
5.8948e-315 0
0
6 74LS95
110 1217 254 0 12 25
0 18 7 7 14 5 6 6 10 8
9 12 13
0
0 0 4336 0
6 74LS95
-21 -51 21 -43
3 U10
-11 -52 10 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7444 0 0
2
5.8948e-315 0
0
6 74LS95
110 1058 254 0 12 25
0 18 7 7 2 2 6 6 6 10
11 36 37
0
0 0 4336 0
6 74LS95
-21 -51 21 -43
2 U9
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 6 9 8 5 4 3 2 1 10
11 12 13 6 9 8 5 4 3 2
1 10 11 12 13 0
65 0 0 512 1 0 0 0
1 U
8503 0 0
2
5.8948e-315 0
0
2 +V
167 84 437 0 1 3
0 19
0
0 0 53744 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3440 0 0
2
40346.6 0
0
10 2-In NAND~
219 764 249 0 3 22
0 16 14 26
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 8 0
1 U
3927 0 0
2
40346.6 1
0
10 2-In NAND~
219 765 337 0 3 22
0 16 24 25
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 6 0
1 U
6639 0 0
2
40346.6 2
0
10 2-In NAND~
219 574 229 0 3 22
0 23 22 21
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 5 0
1 U
4497 0 0
2
40346.6 3
0
10 2-In NAND~
219 523 202 0 3 22
0 14 20 23
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 4 7 0
1 U
8698 0 0
2
40346.6 4
0
10 2-In NAND~
219 523 258 0 3 22
0 17 5 22
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 3 7 0
1 U
5654 0 0
2
40346.6 5
0
10 2-In NAND~
219 333 249 0 3 22
0 28 20 27
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 82
65 0 0 0 4 2 7 0
1 U
5435 0 0
2
40346.6 6
0
10 2-In NAND~
219 124 153 0 3 22
0 31 30 29
0
0 0 112 512
6 74LS00
-14 -24 28 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 26
65 0 0 0 4 1 7 0
1 U
9317 0 0
2
40346.6 7
0
6 JK RN~
219 651 266 0 6 22
0 21 18 17 19 28 16
0
0 0 4464 0
2 01
-8 -42 6 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 1 3 0
1 U
7781 0 0
2
5.8948e-315 0
0
10 3-In NAND~
219 194 174 0 4 22
0 14 16 17 30
0
0 0 112 180
6 74LS10
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 4 0
1 U
7156 0 0
2
5.8948e-315 5.26354e-315
0
10 3-In NAND~
219 195 133 0 4 22
0 24 28 20 31
0
0 0 112 180
6 74LS10
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 118
65 0 0 0 3 1 4 0
1 U
7558 0 0
2
5.8948e-315 5.30499e-315
0
7 Pulser~
4 83 372 0 10 12
0 38 39 18 40 0 0 20 20 13
8
0
0 0 4144 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7486 0 0
2
40346.6 8
0
14 Logic Display~
6 605 60 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5754 0 0
2
40346.6 9
0
14 Logic Display~
6 560 60 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
951 0 0
2
40346.6 10
0
14 Logic Display~
6 514 60 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5582 0 0
2
40346.6 11
0
14 Logic Display~
6 467 60 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3966 0 0
2
40346.6 12
0
6 JK RN~
219 860 266 0 6 22
0 26 18 25 19 20 17
0
0 0 4464 0
2 00
-8 -42 6 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
65 0 0 0 2 2 2 0
1 U
7978 0 0
2
5.8948e-315 5.32571e-315
0
6 JK RN~
219 417 266 0 6 22
0 27 18 19 19 24 14
0
0 0 4464 0
2 02
-8 -42 6 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 20729136
65 0 0 0 2 2 1 0
1 U
7307 0 0
2
5.8948e-315 5.34643e-315
0
6 JK RN~
219 205 266 0 6 22
0 29 18 19 19 41 5
0
0 0 4464 0
2 03
-8 -42 6 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 20730052
65 0 0 512 2 1 1 0
1 U
441 0 0
2
5.8948e-315 5.3568e-315
0
73
11 1 3 0 0 8320 0 13 6 0 0 7
1407 282
1420 282
1420 439
1284 439
1284 487
1296 487
1296 486
12 1 4 0 0 8320 0 13 5 0 0 6
1407 291
1407 430
1265 430
1265 487
1275 487
1275 486
5 0 5 0 0 12416 0 14 0 0 59 4
1185 263
1167 263
1167 83
467 83
8 0 6 0 0 4096 0 15 0 0 14 2
1026 290
1002 290
3 0 7 0 0 4096 0 13 0 0 6 2
1337 246
1286 246
0 2 7 0 0 8192 0 0 13 31 0 4
1132 405
1286 405
1286 237
1337 237
1 0 8 0 0 20608 0 7 0 0 22 6
1254 486
1254 487
1243 487
1243 423
1274 423
1274 291
10 1 9 0 0 8320 0 14 8 0 0 6
1249 272
1267 272
1267 417
1221 417
1221 487
1232 487
1 0 10 0 0 16512 0 11 0 0 21 5
1137 487
1126 487
1126 417
1112 417
1112 263
1 10 11 0 0 8320 0 12 15 0 0 4
1114 487
1101 487
1101 272
1090 272
11 1 12 0 0 8320 0 14 9 0 0 6
1249 281
1258 281
1258 387
1170 387
1170 487
1181 487
12 1 13 0 0 4224 0 14 10 0 0 5
1249 290
1249 396
1148 396
1148 487
1159 487
7 0 6 0 0 0 0 15 0 0 14 2
1026 281
1002 281
6 0 6 0 0 8192 0 15 0 0 26 3
1026 272
1002 272
1002 327
7 0 6 0 0 0 0 14 0 0 16 2
1185 281
1167 281
6 0 6 0 0 0 0 14 0 0 26 3
1185 272
1167 272
1167 327
5 0 2 0 0 4096 0 15 0 0 18 2
1026 263
1016 263
4 0 2 0 0 8192 0 15 0 0 25 3
1026 254
1016 254
1016 344
4 0 14 0 0 12416 0 14 0 0 58 4
1185 254
1177 254
1177 93
514 93
9 1 15 0 0 4224 0 13 4 0 0 2
1407 264
1407 136
8 9 10 0 0 0 0 14 15 0 0 4
1185 290
1121 290
1121 263
1090 263
8 9 8 0 0 0 0 13 14 0 0 4
1343 291
1274 291
1274 263
1249 263
7 0 16 0 0 12416 0 13 0 0 57 4
1343 282
1328 282
1328 103
560 103
6 0 17 0 0 12416 0 13 0 0 56 4
1343 273
1317 273
1317 114
605 114
1 5 2 0 0 4224 0 2 13 0 0 4
939 344
1307 344
1307 264
1343 264
4 1 6 0 0 12416 0 13 1 0 0 4
1343 255
1297 255
1297 327
940 327
1 0 18 0 0 8192 0 13 0 0 28 3
1343 228
1343 177
1185 177
1 0 18 0 0 8320 0 14 0 0 29 3
1185 227
1185 177
1026 177
1 0 18 0 0 12288 0 15 0 0 40 5
1026 227
1026 177
913 177
913 363
824 363
3 0 7 0 0 0 0 14 0 0 31 2
1179 245
1132 245
2 0 7 0 0 8320 0 14 0 0 33 4
1179 236
1132 236
1132 405
989 405
3 0 7 0 0 0 0 15 0 0 33 2
1020 245
989 245
2 3 7 0 0 0 0 15 3 0 0 4
1020 236
989 236
989 405
964 405
3 0 19 0 0 4096 0 33 0 0 38 3
393 267
393 306
417 306
3 0 19 0 0 0 0 34 0 0 39 3
181 267
181 306
205 306
0 4 19 0 0 4096 0 0 32 37 0 3
651 446
860 446
860 297
4 0 19 0 0 8320 0 24 0 0 38 3
651 297
651 446
417 446
4 0 19 0 0 0 0 33 0 0 39 3
417 297
417 446
205 446
1 4 19 0 0 0 0 16 34 0 0 3
84 446
205 446
205 297
0 2 18 0 0 4096 0 0 32 41 0 4
605 363
824 363
824 258
829 258
0 2 18 0 0 4224 0 0 24 42 0 4
386 363
606 363
606 258
620 258
0 2 18 0 0 0 0 0 33 43 0 3
174 363
386 363
386 258
2 3 18 0 0 0 0 34 27 0 0 3
174 258
174 363
107 363
1 0 17 0 0 0 0 21 0 0 69 3
499 249
488 249
488 165
2 0 20 0 0 4096 0 20 0 0 68 2
499 211
499 124
3 1 21 0 0 12416 0 19 24 0 0 4
601 229
606 229
606 249
627 249
6 2 5 0 0 0 0 34 21 0 0 6
229 249
262 249
262 323
487 323
487 267
499 267
1 0 14 0 0 0 0 20 0 0 73 2
499 193
441 193
3 2 22 0 0 4224 0 21 19 0 0 2
550 258
550 238
3 1 23 0 0 4224 0 20 19 0 0 2
550 202
550 220
2 6 14 0 0 0 0 17 33 0 0 6
740 258
702 258
702 297
470 297
470 249
441 249
1 0 16 0 0 0 0 17 0 0 54 4
740 240
726 240
726 249
690 249
2 5 24 0 0 12288 0 18 33 0 0 6
741 346
678 346
678 311
461 311
461 267
447 267
1 6 16 0 0 0 0 18 24 0 0 4
741 328
690 328
690 249
675 249
3 0 17 0 0 0 0 24 0 0 69 3
627 267
617 267
617 165
1 0 17 0 0 0 0 28 0 0 69 2
605 78
605 165
1 0 16 0 0 0 0 29 0 0 71 2
560 78
560 174
0 1 14 0 0 0 0 0 30 73 0 4
422 183
422 100
514 100
514 78
6 1 5 0 0 0 0 34 31 0 0 4
229 249
229 90
467 90
467 78
3 3 25 0 0 8320 0 18 32 0 0 4
792 337
793 337
793 267
836 267
3 1 26 0 0 4224 0 17 32 0 0 2
791 249
836 249
1 3 27 0 0 4224 0 33 22 0 0 2
393 249
360 249
0 2 20 0 0 4096 0 0 22 68 0 3
278 124
278 258
309 258
0 1 28 0 0 4096 0 0 22 70 0 3
290 133
290 240
309 240
3 1 29 0 0 8320 0 23 34 0 0 4
99 153
98 153
98 249
181 249
4 2 30 0 0 8320 0 25 23 0 0 4
167 174
158 174
158 162
150 162
4 1 31 0 0 8320 0 26 23 0 0 4
168 133
158 133
158 144
150 144
5 3 20 0 0 8320 0 32 26 0 0 3
890 267
890 124
219 124
6 3 17 0 0 0 0 32 25 0 0 3
884 249
884 165
218 165
5 2 28 0 0 8320 0 24 26 0 0 3
681 267
681 133
219 133
6 2 16 0 0 0 0 24 25 0 0 3
675 249
675 174
218 174
5 1 24 0 0 8320 0 33 26 0 0 3
447 267
447 142
219 142
6 1 14 0 0 0 0 33 25 0 0 3
441 249
441 183
218 183
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
